/* Hint in 1-bit bitwise-NOT(~) and logical-NOT(!) operators are the same */
module inverter(input in, 
                output out);

    assign out = ~in;
    
endmodule
